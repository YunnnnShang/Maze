----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 09/21/2023 01:04:23 PM
-- Design Name: 
-- Module Name: success - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity success is
    Port ( resetn : in STD_LOGIC;
           clk25 : in STD_LOGIC;
           F_End: in boolean;
           HC : in integer range 1 to 800;
           VC : in integer range 1 to 525;
           pixel_data_from_rom : out  std_logic_vector (11 downto 0);
           address: in integer range 0 to 19199;
           pixel_pkq: out  std_logic_vector (11 downto 0)
           );
end success;

architecture Behavioral of success is
 type image_array is array (0 to 19199) of std_logic_vector(11 downto 0);
 type image_pkq is array (0 to 323) of std_logic_vector(11 downto 0);
constant pkq: image_pkq := (
x"0FF", x"0FF", x"0FF", x"0BB", x"055", x"0DD", x"0FF", x"0FF", x"0FF", x"0FF", x"0FF", x"0FF", x"0FF", x"0FF", x"0FF", x"0FF", x"0FF", x"0FF", 
x"0FF", x"0FF", x"0FF", x"0FF", x"033", x"041", x"0FC", x"0FF", x"0FF", x"0FF", x"0FF", x"0FF", x"0FF", x"0FF", x"0FF", x"0FF", x"0FF", x"0FF", 
x"0FF", x"0FF", x"0FF", x"0FF", x"0BC", x"071", x"0E4", x"0FD", x"0FF", x"0FF", x"0FF", x"0FF", x"0FF", x"0FF", x"0FF", x"0FF", x"0FF", x"0FF", 
x"0ED", x"0FF", x"0FF", x"0FF", x"0FF", x"0D9", x"0D1", x"0E5", x"0FE", x"0FF", x"0FF", x"0FF", x"0FF", x"0FE", x"0FB", x"0C8", x"033", x"077", 
x"0EA", x"0EC", x"0FF", x"0FF", x"0FF", x"0FF", x"0D9", x"0D2", x"0D5", x"0E6", x"0E7", x"0EB", x"0E9", x"0D3", x"0E2", x"093", x"088", x"0FF", 
x"0D5", x"0E6", x"0E7", x"0FC", x"0FF", x"0FF", x"0FE", x"0A4", x"0D1", x"0E1", x"0E3", x"0E8", x"0E9", x"0D6", x"0EB", x"0FE", x"0FF", x"0FF", 
x"0D2", x"0D2", x"0D1", x"0D2", x"0EA", x"0FF", x"0DB", x"0C1", x"0D2", x"074", x"0B2", x"0E3", x"0D5", x"0B9", x"0FF", x"0FF", x"0FF", x"0FF", 
x"0D3", x"0E1", x"0D2", x"0D1", x"0D1", x"0E8", x"0D8", x"0A1", x"092", x"093", x"0C2", x"0D2", x"0B2", x"0A5", x"0FF", x"0FF", x"0FF", x"0FF", 
x"0D3", x"0E1", x"0E2", x"0E2", x"0D2", x"0B2", x"0B2", x"092", x"052", x"0C2", x"0E2", x"0D2", x"0E2", x"0B3", x"0EE", x"0FF", x"0FF", x"0FF", 
x"0D8", x"0D3", x"0D2", x"0C2", x"0B2", x"092", x"0B2", x"0B2", x"0B2", x"0B2", x"0C2", x"0D2", x"0D2", x"0D9", x"0FF", x"0FF", x"0FF", x"0FF", 
x"0FF", x"0FF", x"0EC", x"0B3", x"0A2", x"073", x"0A2", x"0C2", x"0C2", x"0C2", x"0C2", x"0D2", x"0D3", x"0FE", x"0FF", x"0FF", x"0FF", x"0FF", 
x"0FF", x"0FF", x"0DA", x"0A2", x"0A6", x"085", x"091", x"0C2", x"0E4", x"0D3", x"0E2", x"0D2", x"0E4", x"0FD", x"0FF", x"0FF", x"0FF", x"0FF", 
x"0FF", x"0FF", x"0FE", x"0C9", x"073", x"093", x"0B2", x"0A2", x"0D3", x"0D3", x"0D2", x"0C2", x"0E5", x"0FE", x"0FF", x"0FF", x"0FF", x"0FF", 
x"0FF", x"0FF", x"0FF", x"0A9", x"043", x"062", x"0C2", x"0D2", x"0B2", x"0D2", x"0D2", x"0C2", x"0D4", x"0FF", x"0FF", x"0FF", x"0FF", x"0FF", 
x"0FF", x"0FF", x"0FF", x"0FF", x"076", x"081", x"0D2", x"0E2", x"0D2", x"0D2", x"0E2", x"0D2", x"0D2", x"0FD", x"0FF", x"0FF", x"0FF", x"0FF", 
x"0FF", x"0FF", x"0FF", x"0FF", x"0FF", x"0A5", x"0B1", x"0D2", x"0D2", x"0D2", x"0D1", x"0D2", x"0D2", x"0FC", x"0FF", x"0FF", x"0FF", x"0FF", 
x"0FF", x"0FF", x"0FF", x"0FF", x"0FF", x"0ED", x"094", x"0A2", x"0B2", x"0B4", x"0B4", x"0A2", x"0B4", x"0FF", x"0FF", x"0FF", x"0FF", x"0FF", 
x"0FF", x"0FF", x"0FF", x"0FF", x"0FF", x"0FF", x"0DB", x"0A6", x"0EE", x"0FF", x"0FF", x"0ED", x"0DB", x"0FF", x"0FF", x"0FF", x"0FF", x"0FF"
);      
        
        
        
        
        constant image_data: image_array := (x"01C", x"01C", x"01D", x"01D", x"01D", x"01D", x"01D", x"01D", x"01C", x"01C", x"01C", x"01D", x"01D", x"01D", x"01D", x"01C", x"01C", x"01C", x"01D", x"01D", x"01D", x"01D", x"01C", x"01D", x"01D", x"01D", x"01D", x"01D", x"01D", x"01D", x"01D", x"01D", x"01D", x"01D", x"01C", x"01C", x"01D", x"01D", x"01C", x"01D", x"01D", x"01D", x"01D", x"01D", x"01D", x"01C", x"01C", x"01D", x"01D", x"01D", x"01D", x"01D", x"01D", x"01D", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01D", x"01D", x"01D", x"01D", x"01D", x"01D", x"01D", x"01D", x"01D", x"01D", x"01D", x"01D", x"01D", x"01D", x"01D", x"01D", x"01D", x"01C", x"01C", x"01D", x"01D", x"01D", x"01C", x"01C", x"01D", x"01D", x"01C", x"01D", x"01C", x"01C", x"01C", x"01D", x"01D", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01D", x"01D", x"01D", x"01C", x"01C", x"01C", x"01C", x"01C", x"01D", x"01D", x"01D", x"01D", x"01D", x"01D", x"01C", x"01D", x"01D", x"01C", x"01C", x"01C", x"01C", 
x"01C", x"01C", x"01D", x"01D", x"01D", x"01D", x"01D", x"01D", x"01D", x"01C", x"01C", x"01D", x"01D", x"01D", x"01D", x"01C", x"01D", x"01D", x"01C", x"01D", x"01D", x"01D", x"01C", x"01C", x"01C", x"01C", x"01C", x"01D", x"01D", x"01D", x"01D", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01D", x"01C", x"01D", x"01D", x"01D", x"01D", x"01D", x"01C", x"01C", x"01C", x"01D", x"01D", x"01D", x"01D", x"01D", x"01D", x"01D", x"01C", x"01C", x"01C", x"01C", x"01C", x"01D", x"01D", x"01D", x"01D", x"01D", x"01D", x"01D", x"01D", x"01D", x"01D", x"01D", x"01C", x"01D", x"01D", x"01D", x"01D", x"01C", x"01C", x"01C", x"01C", x"01D", x"01D", x"01D", x"01C", x"01C", x"01C", x"01C", x"01C", x"01D", x"01C", x"01C", x"01C", x"01D", x"01D", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01D", x"01D", x"01D", x"01C", x"01C", x"01C", x"01C", x"01C", x"01D", x"01D", x"01D", x"01D", x"01D", x"01D", x"01D", x"01D", x"01C", x"01C", x"01C", x"01C", x"01C", 
x"01C", x"01C", x"01C", x"01D", x"01D", x"01D", x"01D", x"01D", x"01D", x"01D", x"01C", x"01C", x"01D", x"01D", x"01C", x"01C", x"01C", x"01C", x"01C", x"01D", x"01D", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01D", x"01D", x"01D", x"01D", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01D", x"01D", x"01D", x"01C", x"01C", x"01C", x"01C", x"01C", x"01D", x"01D", x"01D", x"01D", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01D", x"01D", x"01D", x"01D", x"01D", x"01D", x"01C", x"01C", x"01C", x"01D", x"01D", x"01D", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01D", x"01D", x"01D", x"01C", x"01C", x"01C", x"01C", x"01C", x"01D", x"01D", x"01D", x"01D", x"01C", x"01D", x"01D", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", 
x"01C", x"01C", x"01C", x"01C", x"01D", x"01C", x"01C", x"01D", x"01D", x"01D", x"01C", x"01C", x"01D", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01D", x"01C", x"01D", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01D", x"01C", x"01C", x"01C", x"01C", x"01C", x"01D", x"01D", x"01D", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01D", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01D", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01D", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01D", x"01C", x"01C", x"01D", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", 
x"01C", x"01C", x"01C", x"01C", x"01D", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", 
x"01C", x"01C", x"01C", x"01C", x"01D", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", 
x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01B", x"01B", 
x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01B", x"01B", x"01B", 
x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01B", x"01B", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01B", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01B", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01B", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01B", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01B", x"01B", x"01B", 
x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01B", x"01C", x"01B", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01B", x"01B", x"01B", x"01C", x"01C", x"01C", x"01B", x"01C", x"01C", x"01B", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01B", x"01C", x"01B", x"01C", x"01C", x"01B", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01B", x"01B", x"01B", x"01B", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01B", x"01B", x"01B", x"01B", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01B", x"01B", x"01B", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01B", x"01B", x"01B", x"01B", 
x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01B", x"01C", x"01C", x"01C", x"01B", x"01B", x"01B", x"01B", x"01C", x"01C", x"01C", x"01C", x"01C", x"01B", x"01B", x"01B", x"01B", x"01C", x"01C", x"01B", x"01B", x"01B", x"01C", x"01B", x"01C", x"01C", x"01C", x"01B", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01C", x"01B", x"01B", x"01C", x"01C", x"01C", x"01B", x"01B", x"01B", x"01B", x"01B", x"01C", x"01C", x"01C", x"01C", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01C", x"01C", x"01B", x"01C", x"01C", x"01C", x"01B", x"01B", x"01B", x"01B", x"01B", x"01C", x"01C", x"01C", x"01C", x"01C", x"01B", x"01C", x"01C", x"01B", x"01C", x"01B", x"01B", x"01B", x"01C", x"01B", x"01B", x"01B", x"01B", 
x"01C", x"01C", x"01B", x"01C", x"01B", x"01C", x"01C", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01C", x"01B", x"01B", x"01B", x"01B", x"01B", x"01C", x"01C", x"01B", x"01C", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01C", x"01B", x"01B", x"01B", x"01B", x"01B", x"01C", x"01B", x"01C", x"01C", x"01C", x"01C", x"01B", x"01B", x"01C", x"01C", x"01C", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01C", x"01C", x"01B", x"01C", x"01B", x"01B", x"01B", x"01C", x"01C", x"01B", x"01B", x"01C", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01C", x"01C", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01C", x"01C", x"01B", x"01B", x"01B", x"01B", x"01B", x"01C", x"01C", x"01C", x"01C", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", 
x"01B", x"01B", x"01B", x"01C", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01C", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01C", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01C", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01C", x"01C", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", 
x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", 
x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", 
x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"00B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", 
x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", 
x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"00B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"00B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"00B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"00B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"00B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", 
x"00B", x"00B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"00B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"00B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"00B", x"01B", x"01B", x"00B", x"01B", x"00B", x"01B", x"01B", x"01B", x"00B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"00B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"00B", x"00B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"00B", x"00B", x"01B", x"01B", x"01B", x"01B", x"00B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", 
x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"00B", x"01B", x"01B", x"01B", x"01B", x"01B", x"00B", x"01B", x"00B", x"01B", x"01B", x"00B", x"00B", x"01B", x"01B", x"01B", x"01B", x"00B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"00B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"00B", x"01B", x"01B", x"00B", x"01B", x"00B", x"01B", x"01B", x"01B", x"00B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"00B", x"00B", x"01B", x"00B", x"00B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"00B", x"01B", x"01B", x"00B", x"00B", x"01B", x"01B", x"01B", x"01B", x"00B", x"00B", x"01B", x"01B", x"01B", x"01B", x"00B", x"00B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"00B", x"00B", x"01B", 
x"01B", x"01B", x"01B", x"01B", x"00B", x"00B", x"00B", x"01B", x"00B", x"00B", x"01B", x"00B", x"00B", x"01B", x"00B", x"00B", x"01B", x"01B", x"00B", x"00B", x"01B", x"01B", x"01B", x"00B", x"00B", x"01B", x"01B", x"01B", x"00B", x"01B", x"01B", x"00B", x"00B", x"01B", x"00B", x"01B", x"01B", x"00B", x"01B", x"01B", x"01B", x"01B", x"00B", x"00B", x"00B", x"00B", x"01B", x"01B", x"01B", x"01B", x"00B", x"00B", x"00B", x"01B", x"01B", x"00B", x"01B", x"00B", x"01B", x"01B", x"01B", x"00B", x"01B", x"01B", x"00B", x"00B", x"01B", x"01B", x"01B", x"00B", x"00B", x"01B", x"00B", x"00B", x"00B", x"00B", x"00B", x"01B", x"01B", x"01B", x"01B", x"01B", x"00B", x"01B", x"00B", x"01B", x"01B", x"01B", x"01B", x"00B", x"00B", x"00B", x"01B", x"01B", x"01B", x"01B", x"00B", x"01B", x"01B", x"01B", x"00B", x"01B", x"00B", x"01B", x"00A", x"00B", x"00B", x"00B", x"01B", x"00B", x"00B", x"00B", x"01B", x"00B", x"01B", x"01B", x"01B", x"01B", x"00A", x"01B", 
x"01B", x"01B", x"01B", x"01B", x"00B", x"00B", x"00B", x"00B", x"00B", x"00B", x"00B", x"00B", x"00B", x"01B", x"00B", x"00B", x"01B", x"01B", x"01B", x"00B", x"00B", x"00B", x"00B", x"00B", x"00B", x"01B", x"01B", x"01B", x"00B", x"01B", x"01B", x"00B", x"00B", x"00B", x"00B", x"00B", x"00B", x"01B", x"01B", x"01B", x"01B", x"01B", x"00B", x"00B", x"00B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"00B", x"00B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"00B", x"01B", x"01B", x"01B", x"01B", x"01B", x"00B", x"01B", x"00B", x"00B", x"00B", x"00B", x"00B", x"00B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"00B", x"00B", x"00B", x"00B", x"01B", x"00B", x"00B", x"01B", x"01B", x"01B", x"01B", x"00B", x"01B", x"00B", x"01B", x"00B", x"01B", x"00B", x"01B", x"00B", x"00B", x"00B", x"00B", x"01B", x"00B", x"01B", x"00B", x"00B", x"00B", x"00B", x"01B", x"01B", x"01B", x"01B", x"01B", 
x"01B", x"01B", x"01B", x"00B", x"00B", x"00B", x"00B", x"00B", x"00B", x"00B", x"00B", x"00B", x"00B", x"01B", x"01B", x"00B", x"00B", x"01B", x"01B", x"00B", x"00B", x"00B", x"00B", x"00B", x"01B", x"00B", x"01B", x"01B", x"00B", x"01B", x"01B", x"00B", x"00B", x"00B", x"00B", x"00B", x"00B", x"01B", x"01B", x"00B", x"00B", x"00B", x"00B", x"00B", x"01B", x"01B", x"01B", x"00B", x"01B", x"00B", x"01B", x"01B", x"00B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"00B", x"01B", x"01B", x"01B", x"00B", x"00B", x"00B", x"01B", x"00B", x"01B", x"00B", x"01B", x"00B", x"01B", x"00B", x"00B", x"00B", x"00B", x"00B", x"00B", x"01B", x"01B", x"00B", x"01B", x"01B", x"01B", x"00B", x"00B", x"00B", x"00B", x"00B", x"00B", x"00B", x"00B", x"00B", x"01B", x"01B", x"00B", x"01B", x"00B", x"00B", x"00B", x"00B", x"00B", x"01B", x"00B", x"00B", x"01B", x"00B", x"01B", x"00B", x"00B", x"00B", x"00B", x"01B", x"00B", x"01B", x"01B", x"01B", x"00B", x"01A", 
x"01B", x"01B", x"01B", x"00B", x"00A", x"00B", x"00B", x"00B", x"00B", x"00B", x"00B", x"01B", x"01B", x"00B", x"00B", x"00B", x"01B", x"00B", x"01B", x"00B", x"00B", x"00B", x"01B", x"01B", x"01B", x"00B", x"00B", x"01B", x"00B", x"00B", x"00B", x"00B", x"00B", x"00B", x"01B", x"01B", x"01B", x"00B", x"01B", x"00B", x"00A", x"00B", x"00B", x"00B", x"00B", x"01B", x"00B", x"00B", x"01B", x"00B", x"01B", x"01B", x"00B", x"01B", x"01B", x"00B", x"00B", x"00B", x"01B", x"00B", x"00B", x"01B", x"01B", x"00A", x"00A", x"00A", x"00B", x"00B", x"00A", x"00A", x"00B", x"00A", x"01B", x"01B", x"00B", x"00B", x"00B", x"00B", x"00B", x"01B", x"01B", x"00B", x"00B", x"01B", x"00B", x"00B", x"00B", x"00B", x"00B", x"00B", x"00B", x"00B", x"00B", x"00B", x"00B", x"00B", x"00A", x"01B", x"01B", x"00B", x"00B", x"00B", x"00B", x"01B", x"00B", x"00B", x"00B", x"00B", x"01B", x"00B", x"00B", x"00B", x"00B", x"01B", x"00B", x"00B", x"00B", x"00B", x"00A", x"00A", 
x"00B", x"01B", x"00A", x"00A", x"00A", x"00B", x"00B", x"00A", x"00A", x"00A", x"00A", x"00A", x"00B", x"00A", x"00A", x"00B", x"00B", x"00A", x"00B", x"00A", x"00A", x"00B", x"01B", x"01B", x"01B", x"00B", x"00A", x"00B", x"00B", x"00A", x"00A", x"00B", x"00B", x"00B", x"00B", x"00B", x"01B", x"01A", x"00A", x"00A", x"00A", x"00A", x"00B", x"00B", x"00A", x"00B", x"00A", x"00B", x"01B", x"01B", x"00B", x"01B", x"00B", x"00B", x"00B", x"00B", x"00A", x"00A", x"00A", x"00A", x"00A", x"01A", x"01A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"01A", x"01A", x"00B", x"00B", x"00B", x"00B", x"00B", x"00B", x"00A", x"00B", x"00B", x"00B", x"00B", x"00B", x"00B", x"00B", x"00B", x"00B", x"00B", x"00B", x"00B", x"00B", x"00B", x"00B", x"00B", x"00B", x"00A", x"01A", x"01B", x"00A", x"00A", x"00A", x"00B", x"00B", x"00B", x"00B", x"00A", x"00A", x"00B", x"00A", x"00B", x"00B", x"00B", x"00B", x"00B", x"00B", x"00B", x"01B", x"01A", x"00A", 
x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00B", x"00A", x"01B", x"00A", x"00A", x"00A", x"00A", x"00B", x"00B", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00B", x"00A", x"00A", x"00A", x"00A", x"00B", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00B", x"00B", x"00B", x"00A", x"00A", x"00B", x"00B", x"00A", x"01B", x"01B", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"01A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"01A", x"00A", x"00A", x"00A", x"00B", x"01B", x"00B", x"00A", x"00B", x"00B", x"00B", x"00A", x"00A", x"01B", x"00B", x"00A", x"00A", x"00A", x"00A", x"00B", x"01B", x"00B", x"00A", x"00B", x"00B", x"00A", x"00A", x"01A", x"00A", x"00A", x"00A", x"00B", x"00A", x"00B", x"00A", x"00A", x"00A", x"00A", x"00A", x"00B", x"00B", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"01A", x"00A", 
x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00B", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00B", x"01B", x"00A", x"00A", x"00A", x"00A", x"00A", x"01B", x"01A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00B", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", 
x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"01B", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", 
x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", 
x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", 
x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", 
x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", 
x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", 
x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", 
x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", 
x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", 
x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", 
x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", 
x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", 
x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"01A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", 
x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"009", 
x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"009", x"009", 
x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"009", x"009", 
x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"009", x"009", 
x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"01A", x"00A", x"00A", x"00A", x"00A", x"01A", x"00A", x"00A", x"01A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"01A", x"01A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"009", x"009", x"009", 
x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"01A", x"00A", x"00A", x"00A", x"00A", x"01A", x"00A", x"00A", x"00A", x"01A", x"01A", x"00A", x"00A", x"00A", x"00A", x"01A", x"01A", x"01A", x"00A", x"00A", x"00A", x"00A", x"01A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"01A", x"00A", x"00A", x"01A", x"00A", x"00A", x"01A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"009", x"009", 
x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"009", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"01A", x"00A", x"00A", x"00A", x"00A", x"01A", x"00A", x"01A", x"00A", x"01A", x"01A", x"01A", x"01A", x"01A", x"00A", x"01A", x"01A", x"01A", x"00A", x"00A", x"00A", x"00A", x"01A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"01A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"00A", x"00A", x"01A", x"01A", x"00A", x"01A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"009", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"009", x"009", 
x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"009", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"01A", x"00A", x"00A", x"00A", x"00A", x"00A", x"01A", x"00A", x"00A", x"00A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"00A", x"00A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"01A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"00A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"00A", x"01A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"009", x"00A", x"00A", x"00A", x"00A", x"00A", x"009", x"009", x"009", 
x"009", x"009", x"00A", x"00A", x"009", x"009", x"009", x"00A", x"00A", x"009", x"009", x"00A", x"009", x"009", x"009", x"00A", x"00A", x"009", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"01A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"00A", x"01A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"009", x"009", x"00A", x"00A", x"00A", x"00A", x"009", x"009", x"009", 
x"009", x"00A", x"00A", x"009", x"00A", x"009", x"009", x"00A", x"009", x"00A", x"00A", x"009", x"009", x"009", x"009", x"009", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"00A", x"00A", x"00A", x"00A", x"01A", x"00A", x"00A", x"00A", x"00A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"00A", x"01A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"009", x"00A", x"009", x"009", x"009", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"009", x"009", x"009", 
x"009", x"00A", x"00A", x"009", x"00A", x"00A", x"009", x"00A", x"009", x"00A", x"00A", x"009", x"009", x"009", x"009", x"009", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"009", x"00A", x"00A", x"00A", x"00A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"00A", x"01A", x"01A", x"01A", x"01A", x"00A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"009", x"00A", x"009", x"009", x"009", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"009", x"009", x"009", 
x"00A", x"00A", x"009", x"009", x"00A", x"00A", x"00A", x"009", x"009", x"00A", x"009", x"00A", x"00A", x"009", x"009", x"009", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"00A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"009", x"00A", x"00A", x"009", x"009", x"009", x"009", x"009", x"009", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"009", x"009", x"009", 
x"00A", x"00A", x"009", x"009", x"00A", x"00A", x"00A", x"00A", x"009", x"009", x"009", x"00A", x"00A", x"009", x"009", x"009", x"00A", x"00A", x"009", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01B", x"01A", x"01A", x"01A", x"01B", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"009", x"00A", x"00A", x"009", x"009", x"00A", x"00A", x"009", x"00A", x"00A", x"00A", x"00A", x"00A", x"009", x"00A", x"00A", x"00A", x"00A", x"009", x"009", 
x"00A", x"009", x"009", x"009", x"00A", x"00A", x"009", x"00A", x"00A", x"009", x"009", x"00A", x"00A", x"009", x"00A", x"00A", x"009", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01B", x"01B", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01B", x"01A", x"01A", x"01B", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"009", x"009", x"00A", x"00A", x"00A", x"009", x"00A", x"00A", x"009", x"009", x"00A", x"00A", x"00A", x"00A", x"009", x"009", 
x"00A", x"009", x"009", x"00A", x"00A", x"00A", x"009", x"00A", x"00A", x"009", x"009", x"00A", x"00A", x"009", x"00A", x"00A", x"009", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01B", x"01B", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01B", x"01B", x"01B", x"01B", x"01A", x"01A", x"01A", x"01A", x"01A", x"01B", x"01A", x"01B", x"01B", x"01B", x"01A", x"01B", x"01B", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"009", x"009", x"00A", x"00A", x"00A", x"009", x"009", x"00A", x"009", x"009", x"00A", x"00A", x"00A", x"009", x"009", x"009", 
x"00A", x"00A", x"00A", x"00A", x"00A", x"009", x"009", x"009", x"009", x"009", x"009", x"00A", x"00A", x"00A", x"00A", x"009", x"009", x"00A", x"009", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01A", x"01B", x"01A", x"02B", x"01B", x"02B", x"01B", x"01B", x"01B", x"01B", x"01A", x"01A", x"01B", x"01B", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01B", x"01B", x"01A", x"01B", x"01B", x"02B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"02B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01B", x"01A", x"01A", x"01A", x"01A", x"01A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"009", x"009", x"00A", x"00A", x"009", x"009", x"00A", x"009", x"009", x"009", x"00A", x"00A", x"00A", x"009", x"009", x"009", 
x"00A", x"00A", x"00A", x"00A", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"00A", x"00A", x"00A", x"009", x"009", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02A", x"02A", x"02B", x"02A", x"02B", x"02B", x"01A", x"01A", x"01A", x"01A", x"01A", x"01B", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01B", x"01A", x"01A", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"01B", x"02B", x"02B", x"01B", x"01B", x"01B", x"01A", x"01A", x"01A", x"01A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"009", x"00A", x"009", x"009", x"00A", x"00A", x"009", x"009", x"009", x"009", x"009", x"00A", x"009", x"009", x"009", x"009", x"009", x"009", 
x"00A", x"00A", x"009", x"009", x"009", x"009", x"00A", x"00A", x"009", x"009", x"009", x"009", x"00A", x"009", x"00A", x"00A", x"009", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02A", x"02B", x"02A", x"02B", x"02B", x"02A", x"02A", x"02B", x"02B", x"02B", x"01B", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"01B", x"01A", x"01A", x"01A", x"01A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"009", x"00A", x"00A", x"009", x"00A", x"00A", x"009", x"009", x"009", x"009", x"009", x"00A", x"009", x"009", x"009", x"009", x"009", x"009", 
x"00A", x"009", x"009", x"009", x"009", x"009", x"00A", x"00A", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"01A", x"02A", x"01A", x"01A", x"01B", x"01A", x"01A", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"01B", x"01A", x"01A", x"01A", x"01A", x"01A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"009", x"009", x"009", x"009", x"00A", x"00A", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", 
x"009", x"009", x"009", x"009", x"009", x"009", x"00A", x"00A", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"00A", x"009", x"00A", x"00A", x"00A", x"00A", x"00A", x"01A", x"01A", x"01A", x"01A", x"01A", x"02A", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02A", x"02B", x"02A", x"01A", x"02B", x"02A", x"02A", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"00A", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", 
x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"00A", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"00A", x"00A", x"00A", x"00A", x"00A", x"01A", x"01A", x"01A", x"01A", x"02A", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02A", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02A", x"01A", x"01A", x"01A", x"01A", x"01A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"009", x"009", x"009", x"009", x"009", x"009", x"00A", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", 
x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"00A", x"00A", x"00A", x"00A", x"01A", x"01A", x"01A", x"01A", x"01A", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"02B", x"02B", x"02B", x"02B", x"01A", x"01A", x"01A", x"01A", x"01A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"00A", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", 
x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"00A", x"00A", x"00A", x"01A", x"01A", x"01A", x"01A", x"02B", x"02B", x"02B", x"02B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"02B", x"02B", x"02B", x"02A", x"01A", x"01A", x"01A", x"01A", x"01A", x"00A", x"00A", x"00A", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", 
x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"00A", x"00A", x"009", x"009", x"00A", x"00A", x"00A", x"01A", x"01A", x"01A", x"02B", x"02B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03C", x"03C", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03C", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"02B", x"02B", x"02A", x"01A", x"01A", x"01A", x"01A", x"00A", x"00A", x"00A", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", 
x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"00A", x"00A", x"00A", x"01A", x"01A", x"01A", x"01A", x"02B", x"02B", x"02B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03C", x"03C", x"04C", x"03C", x"03C", x"04C", x"04C", x"03C", x"03C", x"03C", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"02B", x"02B", x"02B", x"02B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"04C", x"04C", x"04C", x"03B", x"04C", x"04C", x"04C", x"03B", x"03C", x"03B", x"04C", x"04C", x"04C", x"04C", x"04C", x"03C", x"03C", x"03B", x"03B", x"03B", x"03B", x"02B", x"01A", x"01A", x"01A", x"01A", x"01A", x"00A", x"00A", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", 
x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"00A", x"00A", x"01A", x"01A", x"01A", x"01A", x"02B", x"02B", x"03B", x"03B", x"03B", x"03C", x"04B", x"03B", x"03B", x"04C", x"04C", x"04C", x"04C", x"04C", x"04C", x"04C", x"04C", x"04C", x"04C", x"04C", x"04C", x"04C", x"04C", x"03C", x"04C", x"03C", x"03B", x"03C", x"03B", x"03B", x"03B", x"02B", x"03B", x"03B", x"03B", x"04B", x"04B", x"04C", x"04C", x"04C", x"04C", x"04C", x"04C", x"04C", x"04C", x"04C", x"04C", x"04C", x"04C", x"04C", x"04C", x"04C", x"04C", x"04C", x"04C", x"04C", x"04C", x"04C", x"03C", x"03C", x"03B", x"03B", x"02B", x"02A", x"01A", x"01A", x"01A", x"01A", x"00A", x"00A", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", 
x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"00A", x"00A", x"01A", x"01A", x"01A", x"01A", x"02B", x"02B", x"03B", x"03C", x"04C", x"04C", x"04C", x"04C", x"04C", x"04C", x"04C", x"04C", x"04C", x"04C", x"05C", x"04C", x"04C", x"04C", x"04C", x"04C", x"04C", x"04C", x"04C", x"04C", x"04C", x"04C", x"04C", x"04C", x"03C", x"03B", x"03B", x"03B", x"03B", x"03B", x"04C", x"04C", x"04C", x"04C", x"04C", x"04C", x"04C", x"04C", x"04C", x"04C", x"04C", x"04C", x"05C", x"05C", x"05C", x"05C", x"05C", x"04C", x"05C", x"05C", x"05C", x"05C", x"04C", x"04C", x"04C", x"04C", x"04C", x"03B", x"03B", x"02A", x"01A", x"01A", x"01A", x"01A", x"00A", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", 
x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"00A", x"01A", x"01A", x"01A", x"02A", x"02B", x"03B", x"03B", x"04C", x"05C", x"05C", x"04C", x"04C", x"05C", x"05C", x"05C", x"04C", x"05C", x"05C", x"05C", x"05C", x"05C", x"05D", x"05C", x"05C", x"05C", x"05C", x"05C", x"04C", x"04C", x"05C", x"05C", x"04C", x"04C", x"03B", x"03C", x"03C", x"03B", x"03C", x"04C", x"05C", x"05C", x"04C", x"04C", x"04C", x"04C", x"05C", x"05C", x"05C", x"05C", x"05C", x"05C", x"05C", x"05C", x"05C", x"05C", x"05C", x"05C", x"05C", x"05C", x"05C", x"05C", x"05C", x"05C", x"05C", x"04C", x"03B", x"03B", x"02A", x"02A", x"01A", x"01A", x"01A", x"00A", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", 
x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"00A", x"00A", x"01A", x"01A", x"01A", x"02A", x"02B", x"03B", x"04C", x"05C", x"05C", x"05C", x"05C", x"05C", x"05C", x"06C", x"05C", x"05C", x"05C", x"06C", x"06C", x"06C", x"06C", x"06C", x"05C", x"05C", x"05C", x"06C", x"06C", x"05C", x"05C", x"05C", x"05C", x"05C", x"04C", x"03B", x"03C", x"03C", x"03C", x"04C", x"05C", x"05C", x"05C", x"05C", x"05C", x"05C", x"05C", x"05C", x"06C", x"06C", x"06C", x"06C", x"06C", x"06C", x"06C", x"06C", x"06C", x"06C", x"06C", x"06C", x"06C", x"06C", x"06C", x"06C", x"06C", x"06C", x"05C", x"04B", x"03B", x"02B", x"02A", x"01A", x"01A", x"01A", x"00A", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", 
x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"00A", x"00A", x"01A", x"01A", x"01A", x"02A", x"02B", x"03B", x"05C", x"08E", x"09E", x"08D", x"06C", x"06C", x"09E", x"0AE", x"08D", x"06C", x"06D", x"09E", x"09E", x"0AE", x"0AE", x"09E", x"07D", x"05C", x"07D", x"09E", x"09E", x"06C", x"05B", x"08D", x"09E", x"08E", x"05C", x"04B", x"03B", x"03B", x"03B", x"04C", x"07D", x"09E", x"09E", x"06C", x"06C", x"06D", x"06C", x"07D", x"09E", x"09E", x"07C", x"08D", x"0AE", x"0AE", x"0AE", x"09E", x"08D", x"07C", x"0AE", x"09E", x"0AE", x"08D", x"06C", x"07D", x"09E", x"09E", x"07C", x"04B", x"03B", x"02B", x"02B", x"01A", x"01A", x"01A", x"00A", x"00A", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", 
x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"00A", x"00A", x"01A", x"01A", x"01A", x"02A", x"02B", x"03B", x"05B", x"0BF", x"0CF", x"0AE", x"06B", x"07D", x"0CF", x"0DF", x"0AE", x"06C", x"07D", x"0BF", x"0CF", x"0DF", x"0DF", x"0CF", x"07C", x"06B", x"09E", x"0CF", x"0CF", x"07C", x"06B", x"0AE", x"0CF", x"0BF", x"06B", x"04B", x"03B", x"03B", x"04B", x"05B", x"0AE", x"0CF", x"0BF", x"07C", x"06C", x"06C", x"06C", x"09E", x"0CF", x"0CF", x"08C", x"0AE", x"0DF", x"0CF", x"0CF", x"0CF", x"09D", x"08C", x"0CF", x"0CF", x"0CF", x"0AE", x"06B", x"09D", x"0CF", x"0CF", x"08D", x"04B", x"03C", x"02B", x"02B", x"02A", x"01A", x"01A", x"01A", x"00A", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", 
x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"00A", x"00A", x"01A", x"01A", x"01A", x"02A", x"02B", x"04B", x"05C", x"0BF", x"0DF", x"0BE", x"06B", x"07D", x"0DF", x"0DF", x"0BD", x"06B", x"08D", x"0CF", x"0DF", x"0DF", x"0DF", x"0DF", x"08C", x"06B", x"0AE", x"0DF", x"0DF", x"08C", x"06B", x"0BF", x"0DF", x"0CF", x"06B", x"04B", x"04B", x"03B", x"04C", x"05C", x"0AF", x"0DF", x"0CF", x"07B", x"07C", x"07C", x"07C", x"0AE", x"0DF", x"0DF", x"08C", x"0AE", x"0DF", x"0DF", x"0DF", x"0DF", x"09D", x"09C", x"0DF", x"0DF", x"0EF", x"0BD", x"07B", x"09D", x"0DF", x"0DF", x"08D", x"04B", x"03C", x"02B", x"02B", x"02A", x"01A", x"01A", x"01A", x"00A", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", 
x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"00A", x"01A", x"01A", x"01A", x"02A", x"02B", x"04C", x"06C", x"0BF", x"0DF", x"0BE", x"07B", x"07D", x"0CF", x"0DF", x"0BD", x"07C", x"0AE", x"0DF", x"0DF", x"0CE", x"0DF", x"0DF", x"0BE", x"08C", x"0AD", x"0DF", x"0DF", x"08C", x"06B", x"0BF", x"0DF", x"0CF", x"06B", x"05B", x"04C", x"04C", x"04C", x"06C", x"0AF", x"0DF", x"0CE", x"08B", x"0AE", x"0BF", x"09D", x"0AE", x"0DF", x"0DF", x"08C", x"0AD", x"0CF", x"0DF", x"0DF", x"0DF", x"09D", x"09C", x"0DF", x"0DF", x"0DF", x"0CE", x"0AD", x"0AD", x"0DF", x"0DF", x"09D", x"05B", x"03B", x"03B", x"02B", x"02A", x"01A", x"01A", x"01A", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", 
x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"00A", x"00A", x"01A", x"01A", x"01A", x"02A", x"03B", x"04C", x"06C", x"0BF", x"0EF", x"0CE", x"07B", x"08D", x"0CF", x"0EF", x"0BD", x"08C", x"0CF", x"0DF", x"0BD", x"08A", x"0AD", x"0DF", x"0DF", x"09C", x"0AD", x"0DF", x"0DF", x"08C", x"07B", x"0BF", x"0EF", x"0CF", x"06B", x"05B", x"04C", x"04C", x"04C", x"06C", x"0BF", x"0DF", x"0DE", x"09B", x"0CF", x"0DF", x"0AD", x"0AD", x"0DF", x"0DF", x"09C", x"07B", x"0AD", x"0DF", x"0DF", x"0AC", x"07B", x"09D", x"0DF", x"0DF", x"0DF", x"0DF", x"0BE", x"0AC", x"0DF", x"0DF", x"09D", x"05B", x"04B", x"03B", x"02B", x"02A", x"01A", x"01A", x"00A", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", 
x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"00A", x"00A", x"01A", x"01A", x"01A", x"02A", x"03B", x"04C", x"06C", x"0BF", x"0EF", x"0CE", x"07B", x"08D", x"0DF", x"0EF", x"0BD", x"09C", x"0DF", x"0EF", x"0BD", x"069", x"09C", x"0DF", x"0DF", x"09C", x"0AD", x"0EF", x"0DF", x"08C", x"07B", x"0BF", x"0EF", x"0CF", x"06B", x"05C", x"04C", x"04C", x"04C", x"06C", x"0BF", x"0EF", x"0DE", x"0AC", x"0DF", x"0EF", x"0BD", x"0BD", x"0EF", x"0DF", x"09D", x"07A", x"09C", x"0EF", x"0DF", x"09B", x"06B", x"0AD", x"0DF", x"0EF", x"0EF", x"0EF", x"0CE", x"0AC", x"0DF", x"0EF", x"09D", x"05B", x"04B", x"03B", x"02B", x"02A", x"01A", x"01A", x"00A", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", 
x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"00A", x"01A", x"01A", x"02A", x"02B", x"03B", x"04C", x"06C", x"0BF", x"0EF", x"0CE", x"08C", x"08D", x"0DF", x"0EF", x"0BD", x"09C", x"0DF", x"0EF", x"0BD", x"08B", x"0AE", x"0DF", x"0DF", x"09C", x"0BD", x"0EF", x"0DF", x"09C", x"07B", x"0BF", x"0EF", x"0CF", x"07B", x"05C", x"04C", x"04C", x"05C", x"06C", x"0BF", x"0EF", x"0DE", x"0AC", x"0DF", x"0DF", x"0BD", x"0BD", x"0EF", x"0DF", x"09D", x"07B", x"0AE", x"0EF", x"0DF", x"09C", x"07C", x"0AD", x"0DF", x"0EF", x"0EF", x"0EF", x"0CE", x"0AC", x"0DF", x"0EF", x"09D", x"05C", x"04C", x"03B", x"02B", x"02A", x"01A", x"01A", x"01A", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", 
x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"00A", x"01A", x"01A", x"01A", x"02B", x"03B", x"04B", x"06C", x"0BF", x"0EF", x"0CE", x"07B", x"08D", x"0DF", x"0EF", x"0BD", x"09C", x"0DF", x"0EF", x"0BD", x"07B", x"0AE", x"0DF", x"0EF", x"0AC", x"0BD", x"0EF", x"0EF", x"09C", x"07B", x"0BF", x"0EF", x"0DF", x"07B", x"05C", x"04C", x"04C", x"05C", x"06C", x"0BF", x"0EF", x"0DE", x"0AB", x"0DF", x"0EF", x"0BD", x"0BC", x"0EF", x"0DF", x"09D", x"07C", x"0AE", x"0EF", x"0DF", x"09C", x"07C", x"0AE", x"0EF", x"0EF", x"0EF", x"0EF", x"0CE", x"0AC", x"0DF", x"0EF", x"09D", x"05B", x"04C", x"03B", x"02B", x"02A", x"01A", x"01A", x"01A", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", 
x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"01A", x"01A", x"01A", x"02B", x"03B", x"04B", x"06C", x"0CF", x"0EF", x"0CE", x"09C", x"0AD", x"0DF", x"0EF", x"0BD", x"09C", x"0DF", x"0EF", x"0BD", x"07B", x"0AE", x"0EF", x"0EF", x"0AC", x"0BD", x"0EF", x"0EF", x"09C", x"07B", x"0BF", x"0EF", x"0DF", x"07B", x"05C", x"04C", x"04C", x"05C", x"06C", x"0BF", x"0EF", x"0DE", x"0BC", x"0DE", x"0EF", x"0CD", x"0CD", x"0EF", x"0DF", x"09D", x"07C", x"0AE", x"0EF", x"0DF", x"09D", x"07D", x"0AE", x"0EF", x"0EF", x"0EF", x"0EF", x"0CE", x"0BD", x"0EF", x"0EF", x"09D", x"05C", x"04C", x"03B", x"02B", x"02A", x"01A", x"01A", x"01A", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", 
x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"01A", x"01A", x"01A", x"02B", x"03B", x"03B", x"05C", x"0AE", x"0DE", x"0DE", x"0CE", x"0CE", x"0DF", x"0CE", x"0AC", x"09C", x"0DF", x"0EF", x"0BD", x"07B", x"0AE", x"0EF", x"0EF", x"0AC", x"0BD", x"0EF", x"0EF", x"09C", x"07C", x"0CF", x"0EF", x"0DF", x"07B", x"05C", x"04C", x"04C", x"05C", x"06C", x"0BF", x"0EF", x"0DE", x"0DE", x"0EF", x"0EF", x"0DE", x"0DE", x"0EF", x"0EF", x"09D", x"07C", x"0AE", x"0EF", x"0EF", x"09D", x"07D", x"0AE", x"0EF", x"0EF", x"0DE", x"0DE", x"0DE", x"0DE", x"0EF", x"0EF", x"09D", x"05C", x"04C", x"03B", x"02B", x"02A", x"01A", x"01A", x"01A", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", 
x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"01A", x"01A", x"01A", x"02A", x"03B", x"04B", x"05C", x"07B", x"0BD", x"0EF", x"0EF", x"0EF", x"0EF", x"0AD", x"07A", x"09D", x"0DF", x"0EF", x"0BD", x"07B", x"0AE", x"0EF", x"0EF", x"0AC", x"0BD", x"0EF", x"0EF", x"09D", x"08C", x"0CF", x"0EF", x"0DF", x"07B", x"05C", x"04C", x"04C", x"05C", x"06C", x"0BF", x"0EF", x"0EF", x"0EF", x"0EF", x"0EF", x"0EF", x"0EF", x"0EF", x"0EF", x"09D", x"07C", x"0AE", x"0EF", x"0EF", x"09D", x"07C", x"0AE", x"0EF", x"0EF", x"0BC", x"0CD", x"0EF", x"0EF", x"0EF", x"0EF", x"0AD", x"06C", x"04C", x"03B", x"02B", x"02A", x"01A", x"01A", x"01A", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", 
x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"00A", x"00A", x"01A", x"01A", x"02A", x"02B", x"03B", x"05C", x"06B", x"0BE", x"0EF", x"0EF", x"0EF", x"0EF", x"0AD", x"07B", x"09D", x"0DF", x"0EF", x"0BD", x"07B", x"0AE", x"0EF", x"0EF", x"0AC", x"0BD", x"0EF", x"0EF", x"09D", x"08C", x"0CF", x"0EF", x"0DF", x"07B", x"05C", x"04C", x"04C", x"05C", x"06C", x"0BF", x"0EF", x"0EF", x"0EF", x"0EF", x"0EF", x"0EF", x"0EF", x"0EF", x"0EF", x"09D", x"07C", x"0AE", x"0EF", x"0EF", x"09C", x"07D", x"0AE", x"0EF", x"0EF", x"0BC", x"0CD", x"0EF", x"0EF", x"0EE", x"0EF", x"0AD", x"05B", x"04B", x"03B", x"02B", x"02A", x"01A", x"01A", x"01A", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", 
x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"00A", x"00A", x"01A", x"01A", x"02A", x"02B", x"03B", x"04B", x"06C", x"09D", x"0CE", x"0EF", x"0EF", x"0CD", x"08C", x"07C", x"09D", x"0DF", x"0EF", x"0BD", x"07B", x"0AE", x"0EF", x"0EF", x"0AC", x"0BD", x"0EF", x"0EF", x"09D", x"08C", x"0CF", x"0EF", x"0DF", x"07B", x"05C", x"04C", x"04C", x"04C", x"06C", x"0BF", x"0EF", x"0EF", x"0EF", x"0EF", x"0EF", x"0EF", x"0EF", x"0EF", x"0EF", x"09D", x"07C", x"0AE", x"0EF", x"0EF", x"09C", x"07C", x"0AE", x"0EF", x"0EF", x"0BD", x"0CE", x"0EF", x"0EE", x"0EF", x"0EF", x"0AD", x"05C", x"04B", x"03B", x"02B", x"02A", x"01A", x"01A", x"01A", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", 
x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"00A", x"01A", x"01A", x"01A", x"02A", x"02B", x"03B", x"04C", x"06C", x"07B", x"0AD", x"0EF", x"0EF", x"0AC", x"07B", x"07C", x"09D", x"0DF", x"0EF", x"0BD", x"07B", x"0AE", x"0EF", x"0EF", x"0AC", x"0BD", x"0EF", x"0EF", x"0AD", x"08C", x"0CF", x"0EF", x"0DF", x"07B", x"05C", x"04C", x"04C", x"04C", x"06C", x"0BF", x"0EF", x"0EF", x"0EF", x"0EF", x"0EF", x"0EF", x"0EF", x"0EF", x"0EF", x"09D", x"07C", x"0AE", x"0EF", x"0EF", x"0AC", x"07C", x"0AE", x"0EF", x"0EF", x"0BD", x"0CE", x"0EF", x"0EE", x"0EF", x"0EF", x"0AD", x"05C", x"04C", x"03B", x"02B", x"02A", x"01A", x"01A", x"01A", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", 
x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"00A", x"01A", x"01A", x"01A", x"02B", x"02B", x"03B", x"04C", x"05C", x"06B", x"0AD", x"0EF", x"0EF", x"09B", x"07B", x"06C", x"09D", x"0DF", x"0EF", x"0BD", x"08B", x"0AE", x"0EF", x"0EF", x"0AC", x"0BD", x"0EF", x"0EF", x"0AD", x"08C", x"0CF", x"0EF", x"0DF", x"07B", x"05C", x"04C", x"04C", x"04C", x"06C", x"0BF", x"0EF", x"0EF", x"0EF", x"0EF", x"0EF", x"0EF", x"0EF", x"0EF", x"0EF", x"09D", x"07C", x"0AE", x"0EF", x"0EF", x"0AC", x"07D", x"0AE", x"0EF", x"0EF", x"0BD", x"0CE", x"0EF", x"0EF", x"0EF", x"0EF", x"09D", x"05C", x"04C", x"03B", x"02B", x"02A", x"01A", x"01A", x"00A", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", 
x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"01A", x"01A", x"01A", x"02B", x"03B", x"03B", x"05C", x"06C", x"0BE", x"0EF", x"0EF", x"09C", x"07C", x"06C", x"09D", x"0DF", x"0EF", x"0BD", x"08B", x"0BE", x"0EF", x"0EF", x"0AC", x"0BD", x"0EF", x"0EF", x"0AC", x"08B", x"0CF", x"0EF", x"0DF", x"07B", x"05C", x"04C", x"04C", x"04C", x"06C", x"09D", x"0CD", x"0EF", x"0EF", x"0CD", x"0BC", x"0DE", x"0EF", x"0EE", x"0BD", x"08C", x"07C", x"0AE", x"0EF", x"0EF", x"0AC", x"07C", x"0AE", x"0EF", x"0EF", x"0BD", x"0AD", x"0CE", x"0EF", x"0EF", x"0EF", x"0AD", x"05C", x"04C", x"03B", x"02B", x"02A", x"01A", x"01A", x"00A", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", 
x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"019", x"01A", x"01A", x"02B", x"02B", x"03C", x"04C", x"06C", x"0AE", x"0EF", x"0EF", x"09C", x"06C", x"06C", x"09D", x"0EF", x"0EF", x"0BD", x"08B", x"0BE", x"0EF", x"0EF", x"0AC", x"0BD", x"0EF", x"0EF", x"0AC", x"09B", x"0CF", x"0EF", x"0DF", x"07B", x"05C", x"04C", x"04C", x"04C", x"05C", x"07C", x"0BD", x"0EF", x"0EF", x"0AC", x"09B", x"0CE", x"0EF", x"0EF", x"08B", x"07C", x"08C", x"0BE", x"0EF", x"0EF", x"0AC", x"08C", x"0AD", x"0EF", x"0EF", x"0BD", x"08C", x"0BE", x"0EF", x"0EF", x"0EF", x"0AD", x"06C", x"04C", x"03B", x"02B", x"02A", x"01A", x"01A", x"00A", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", 
x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"019", x"019", x"01A", x"02B", x"02B", x"03C", x"04C", x"05B", x"0AE", x"0EF", x"0EF", x"09C", x"06B", x"06C", x"08D", x"0DF", x"0EF", x"0CE", x"0AC", x"0CE", x"0EF", x"0DF", x"09C", x"0AD", x"0DF", x"0EF", x"0BD", x"0BD", x"0DF", x"0EF", x"0CF", x"06B", x"05B", x"04C", x"04C", x"04C", x"05C", x"06B", x"0BD", x"0EF", x"0EF", x"0AC", x"08B", x"0CE", x"0EF", x"0DF", x"08B", x"07C", x"09D", x"0CE", x"0EF", x"0EF", x"0BD", x"09D", x"0AD", x"0EF", x"0EF", x"0AD", x"07B", x"0AD", x"0DF", x"0EF", x"0EF", x"0AD", x"06B", x"04B", x"03B", x"02B", x"02A", x"01A", x"01A", x"00A", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", 
x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"00A", x"00A", x"01A", x"019", x"01A", x"02B", x"02B", x"03B", x"04C", x"05B", x"0AE", x"0EF", x"0EF", x"08C", x"06B", x"05C", x"07D", x"0AD", x"0DE", x"0EF", x"0DF", x"0EF", x"0EF", x"0BD", x"08B", x"09C", x"0BD", x"0EF", x"0EF", x"0EF", x"0EF", x"0DE", x"0AC", x"05A", x"04B", x"04B", x"04B", x"04C", x"05C", x"06C", x"0BE", x"0EF", x"0EF", x"0AC", x"08C", x"0CF", x"0EF", x"0DF", x"08B", x"07C", x"0BE", x"0DF", x"0EF", x"0EF", x"0DF", x"0AD", x"0AD", x"0EF", x"0EF", x"0AD", x"07C", x"09D", x"0BD", x"0EF", x"0EF", x"09D", x"05B", x"04B", x"03B", x"02B", x"02A", x"01A", x"01A", x"00A", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", 
x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"00A", x"00A", x"01A", x"01A", x"02A", x"02B", x"03B", x"04C", x"05B", x"0AE", x"0EF", x"0EF", x"09C", x"05B", x"05C", x"06C", x"07B", x"0DF", x"0EF", x"0EF", x"0EF", x"0EF", x"08B", x"06B", x"07B", x"09C", x"0EF", x"0EF", x"0EF", x"0EF", x"0CE", x"069", x"05B", x"04C", x"03B", x"03B", x"04B", x"04C", x"05C", x"0BE", x"0EF", x"0EF", x"09C", x"07B", x"0CF", x"0FF", x"0DF", x"07B", x"07B", x"0BE", x"0EF", x"0EF", x"0EF", x"0EF", x"0AD", x"09C", x"0EF", x"0FF", x"0AC", x"07C", x"07B", x"09C", x"0EF", x"0EF", x"09C", x"05B", x"04B", x"03B", x"02B", x"02A", x"01A", x"019", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", 
x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"00A", x"00A", x"01A", x"01A", x"01A", x"02B", x"03B", x"04B", x"04B", x"09D", x"0CF", x"0DF", x"08B", x"05B", x"05C", x"05C", x"07C", x"0CF", x"0DF", x"0DE", x"0DE", x"0CE", x"07B", x"06C", x"06C", x"09D", x"0CF", x"0DE", x"0DE", x"0DF", x"0BD", x"06A", x"05B", x"04B", x"03B", x"03B", x"03B", x"04C", x"05C", x"0AE", x"0DF", x"0DF", x"08C", x"07B", x"0BE", x"0DF", x"0CE", x"07B", x"06B", x"0AE", x"0DF", x"0DE", x"0DE", x"0DF", x"09D", x"09C", x"0DF", x"0DE", x"09C", x"06B", x"06B", x"09D", x"0DF", x"0DF", x"08C", x"05B", x"03B", x"02B", x"02A", x"01A", x"019", x"019", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", 
x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"00A", x"00A", x"01A", x"01A", x"01A", x"02A", x"02B", x"03B", x"04B", x"07C", x"08C", x"08C", x"06B", x"05B", x"05C", x"05C", x"07C", x"09D", x"09C", x"09C", x"09C", x"09C", x"07C", x"06C", x"06C", x"08D", x"09D", x"09C", x"09C", x"09C", x"08C", x"06B", x"05C", x"04B", x"03B", x"03B", x"03B", x"04C", x"05C", x"07C", x"09C", x"09C", x"06B", x"06C", x"08D", x"09C", x"08C", x"06B", x"06C", x"08D", x"09C", x"09C", x"09C", x"09C", x"07B", x"07C", x"09D", x"09C", x"07B", x"06B", x"06C", x"08D", x"09C", x"09C", x"06B", x"04B", x"03B", x"02B", x"02A", x"01A", x"019", x"019", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", 
x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"01A", x"01A", x"01A", x"02A", x"02B", x"03B", x"04B", x"05B", x"049", x"049", x"04A", x"04C", x"04C", x"05C", x"05C", x"05A", x"04A", x"05A", x"059", x"05A", x"05B", x"05C", x"05C", x"05C", x"05A", x"049", x"059", x"059", x"04A", x"05B", x"04B", x"03B", x"03B", x"03B", x"03B", x"03C", x"04C", x"05B", x"04A", x"049", x"05B", x"06C", x"05B", x"04A", x"04A", x"05B", x"06C", x"05B", x"05A", x"05A", x"05A", x"05A", x"05A", x"06B", x"05A", x"04A", x"05A", x"05C", x"05C", x"06B", x"05A", x"049", x"04A", x"04B", x"03B", x"02B", x"02A", x"01A", x"01A", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", 
x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"019", x"01A", x"01A", x"02A", x"02A", x"02B", x"03B", x"04B", x"05C", x"05C", x"04C", x"04C", x"04C", x"04C", x"05B", x"05C", x"06C", x"06C", x"06C", x"06C", x"05C", x"05C", x"05C", x"05C", x"06C", x"06C", x"06C", x"06C", x"05C", x"05C", x"04B", x"03B", x"03B", x"02B", x"03B", x"03B", x"04C", x"05C", x"05C", x"06C", x"05C", x"05C", x"05C", x"06C", x"06C", x"05C", x"05C", x"05C", x"06C", x"06C", x"06C", x"06C", x"05B", x"05C", x"06C", x"06C", x"05C", x"05C", x"05C", x"05C", x"06C", x"05C", x"04B", x"04B", x"03B", x"02B", x"01A", x"01A", x"01A", x"00A", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", 
x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"01A", x"01A", x"01A", x"02B", x"02B", x"03B", x"04B", x"04C", x"05C", x"04B", x"04B", x"04C", x"04B", x"04B", x"05C", x"05C", x"05C", x"05C", x"05C", x"05C", x"04C", x"04C", x"05C", x"05C", x"05C", x"05C", x"05C", x"04C", x"04C", x"03B", x"03B", x"02B", x"02B", x"02B", x"03B", x"03B", x"04B", x"05B", x"05C", x"05C", x"05C", x"05C", x"05C", x"05C", x"05C", x"04C", x"05C", x"05C", x"05C", x"05C", x"05C", x"05B", x"05C", x"05C", x"05C", x"05C", x"04C", x"04C", x"04C", x"05C", x"04C", x"04B", x"03B", x"02B", x"02B", x"01A", x"01A", x"01A", x"00A", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", 
x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"01A", x"01A", x"01A", x"02A", x"02B", x"03B", x"03B", x"03B", x"04B", x"03B", x"03B", x"03B", x"03B", x"03B", x"04C", x"04C", x"04B", x"04B", x"04B", x"04C", x"04C", x"04B", x"04C", x"04C", x"04C", x"04C", x"04C", x"04B", x"03B", x"03B", x"02B", x"02B", x"02B", x"02B", x"03B", x"03B", x"03B", x"04B", x"04B", x"04B", x"04C", x"04C", x"04C", x"04B", x"04B", x"04B", x"04C", x"04C", x"04C", x"04C", x"04B", x"04B", x"04B", x"04C", x"04C", x"04C", x"04B", x"04B", x"04C", x"04B", x"04B", x"03B", x"03B", x"02A", x"02A", x"01A", x"01A", x"00A", x"00A", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", 
x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"00A", x"01A", x"01A", x"01A", x"01A", x"02B", x"02B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"04B", x"04B", x"04B", x"04C", x"04B", x"04B", x"03B", x"03B", x"04B", x"04C", x"04B", x"04C", x"04B", x"03B", x"03B", x"03B", x"02B", x"02B", x"02B", x"02A", x"02B", x"03B", x"03B", x"03B", x"04B", x"04B", x"03B", x"04B", x"04B", x"04B", x"03B", x"04B", x"04B", x"04C", x"04C", x"04C", x"04B", x"04B", x"04B", x"04C", x"04C", x"04B", x"04B", x"03B", x"03B", x"03C", x"03B", x"03B", x"02B", x"02A", x"02A", x"01A", x"01A", x"00A", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", 
x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"00A", x"00A", x"00A", x"01A", x"01A", x"01A", x"02A", x"02A", x"02A", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"04B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"02B", x"02B", x"02A", x"02A", x"02A", x"02A", x"02B", x"02B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03C", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"02A", x"02A", x"01A", x"01A", x"01A", x"009", x"00A", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", 
x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"00A", x"00A", x"00A", x"01A", x"01A", x"01A", x"01A", x"02A", x"02A", x"02A", x"02B", x"02B", x"02B", x"02B", x"02B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"02B", x"02A", x"02A", x"02A", x"02A", x"02A", x"02A", x"02B", x"02B", x"02B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"02B", x"02A", x"02A", x"02A", x"01A", x"01A", x"00A", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", 
x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"00A", x"00A", x"01A", x"01A", x"01A", x"01A", x"02A", x"02A", x"02A", x"02B", x"02B", x"02B", x"02A", x"02A", x"02B", x"02B", x"03B", x"03B", x"03B", x"02B", x"02B", x"03B", x"03B", x"03B", x"02B", x"02B", x"02B", x"02B", x"02A", x"02A", x"02A", x"02A", x"01A", x"02A", x"02A", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"03B", x"02B", x"02B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"03B", x"02B", x"02B", x"02B", x"02B", x"02A", x"02A", x"02A", x"01A", x"01A", x"01A", x"00A", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", 
x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"00A", x"01A", x"01A", x"01A", x"01A", x"01B", x"02B", x"02A", x"02B", x"02A", x"02A", x"02A", x"02A", x"02A", x"02A", x"02B", x"02B", x"02B", x"02B", x"02A", x"02A", x"02A", x"02B", x"02B", x"02B", x"02B", x"02B", x"02A", x"02A", x"02A", x"01A", x"01A", x"01A", x"01A", x"02A", x"02B", x"02B", x"02B", x"02B", x"02A", x"02A", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02A", x"02A", x"02B", x"02A", x"02B", x"02B", x"02A", x"02A", x"01A", x"01A", x"01A", x"01A", x"00A", x"00A", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", 
x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"00A", x"00A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"02A", x"02A", x"02A", x"02A", x"02A", x"02B", x"02B", x"02B", x"02A", x"02A", x"02A", x"02A", x"02A", x"02B", x"02B", x"02B", x"02A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"02A", x"02A", x"02A", x"02A", x"02A", x"02A", x"02A", x"02A", x"02A", x"02A", x"02B", x"02B", x"02B", x"02B", x"02B", x"02B", x"02A", x"02A", x"02A", x"02B", x"02A", x"02A", x"02B", x"01A", x"01A", x"01A", x"01A", x"01A", x"00A", x"00A", x"00A", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", 
x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"00A", x"00A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"02A", x"02A", x"02A", x"02B", x"02B", x"02A", x"02A", x"02A", x"02A", x"02A", x"02A", x"02A", x"01A", x"02A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"02A", x"02A", x"02A", x"02A", x"02A", x"02B", x"02A", x"02A", x"02A", x"02A", x"02A", x"02A", x"02A", x"02A", x"02A", x"02A", x"02A", x"02A", x"02A", x"02A", x"02A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"00A", x"00A", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", 
x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"00A", x"00A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"02A", x"01A", x"01A", x"02A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"02A", x"02A", x"02A", x"01A", x"01A", x"01A", x"01A", x"01A", x"02A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"019", x"00A", x"00A", x"00A", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", 
x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"00A", x"00A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"00A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"009", x"00A", x"00A", x"00A", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", 
x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"00A", x"00A", x"00A", x"00A", x"01A", x"019", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"00A", x"00A", x"009", x"00A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"00A", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", 
x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"00A", x"01A", x"01A", x"00A", x"009", x"009", x"00A", x"00A", x"00A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"00A", x"00A", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", 
x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"01A", x"01A", x"01A", x"009", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"00A", x"01A", x"01A", x"01A", x"00A", x"00A", x"00A", x"00A", x"00A", x"009", x"009", x"00A", x"00A", x"00A", x"00A", x"00A", x"01A", x"00A", x"01A", x"01A", x"019", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"01A", x"00A", x"00A", x"00A", x"00A", x"00A", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", 
x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"00A", x"00A", x"009", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"009", x"009", x"00A", x"00A", x"01A", x"00A", x"01A", x"00A", x"00A", x"00A", x"009", x"00A", x"00A", x"00A", x"009", x"009", x"009", x"009", x"009", x"00A", x"00A", x"00A", x"00A", x"009", x"00A", x"00A", x"009", x"009", x"00A", x"00A", x"00A", x"01A", x"01A", x"00A", x"00A", x"00A", x"01A", x"01A", x"00A", x"01A", x"01A", x"009", x"009", x"00A", x"00A", x"009", x"009", x"00A", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", 
x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"00A", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"009", x"00A", x"00A", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"009", x"00A", x"00A", x"00A", x"00A", x"009", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"009", x"00A", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", 
x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"00A", x"00A", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", 
x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", 
x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", 
x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", 
x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", 
x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", 
x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", 
x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", 
x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", 
x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", 
x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", 
x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"008", 
x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"008", 
x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", 
x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", 
x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", 
x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", 
x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", 
x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", 
x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", 
x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", 
x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", 
x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", 
x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", 
x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", 
x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", 
x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", 
x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", 
x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", 
x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", 
x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", 
x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", 
x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", 
x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", 
x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", 
x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", 
x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", 
x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", 
x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", 
x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", 
x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", 
x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"00A", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", 
x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"00A", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", 
x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"00A", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"00A", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", 
x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"00A", x"00A", x"009", x"009", x"009", x"00A", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"00A", x"009", x"00A", x"009", x"009", x"00A", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"00A", x"00A", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"00A", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"00A", x"00A", x"009", x"009", x"009", x"009", x"00A", x"009", x"009", x"00A", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", 
x"009", x"009", x"009", x"009", x"009", x"00A", x"00A", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"00A", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"00A", x"00A", x"009", x"009", x"009", x"00A", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"00A", x"009", x"00A", x"009", x"009", x"00A", x"00A", x"00A", x"009", x"009", x"009", x"009", x"009", x"00A", x"00A", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"00A", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"00A", x"00A", x"00A", x"009", x"009", x"00A", x"00A", x"009", x"009", x"00A", x"00A", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", 
x"009", x"009", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"009", x"009", x"009", x"009", x"009", x"009", x"00A", x"00A", x"009", x"00A", x"00A", x"00A", x"00A", x"009", x"00A", x"00A", x"00A", x"00A", x"00A", x"009", x"009", x"009", x"009", x"00A", x"009", x"009", x"009", x"009", x"009", x"00A", x"00A", x"00A", x"009", x"00A", x"00A", x"00A", x"009", x"009", x"009", x"00A", x"00A", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"00A", x"00A", x"00A", x"00A", x"009", x"00A", x"00A", x"00A", x"00A", x"009", x"009", x"009", x"009", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"009", x"009", x"00A", x"00A", x"009", x"00A", x"009", x"009", x"009", x"009", x"009", x"00A", x"00A", x"00A", x"00A", x"009", x"009", x"00A", x"00A", x"00A", x"009", x"00A", x"00A", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"009", x"00A", x"00A", x"009", x"009", x"009", x"009", 
x"009", x"009", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"009", x"009", x"009", x"009", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"009", x"00A", x"00A", x"00A", x"009", x"009", x"00A", x"00A", x"009", x"00A", x"00A", x"00A", x"009", x"009", x"00A", x"00A", x"00A", x"00A", x"00A", x"009", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"009", x"009", x"00A", x"00A", x"00A", x"00A", x"009", x"009", x"009", x"009", x"00A", x"00A", x"00A", x"00A", x"009", x"00A", x"009", x"00A", x"00A", x"009", x"009", x"009", x"009", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"009", x"00A", x"00A", x"009", x"009", x"009", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"009", x"00A", x"00A", x"009", x"009", x"009", x"009", x"009", x"00A", x"009", x"009", x"009", x"009", x"009", x"00A", x"00A", x"00A", x"009", x"009", x"009", 
x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"009", x"009", x"009", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"009", x"009", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"009", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"009", x"009", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"009", x"00A", x"00A", x"00A", x"009", x"009", x"009", x"009", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"009", x"00A", x"00A", x"00A", x"009", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"009", x"009", x"009", x"00A", x"00A", x"00A", x"00A", x"009", x"009", x"009", x"009", x"00A", x"00A", x"00A", x"009", x"009", x"009", 
x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"009", x"009", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"009", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"009", x"00A", x"00A", x"00A", x"009", x"009", x"009", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"009", x"00A", x"00A", x"00A", x"009", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"009", x"009", x"00A", x"00A", x"00A", x"00A", x"009", x"009", x"009", 
x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"009", x"00A", x"00A", x"009", x"009", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"009", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"009", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"009", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"009", x"00A", x"00A", x"00A", x"00A", x"009", x"009", x"009", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"009", x"009", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"00A", x"009", x"00A", x"00A", x"00A", x"009", x"009", x"00A", x"00A", x"00A", x"00A", x"009", x"009", x"009"
);
begin
    process(clk25)
    begin
        if rising_edge (clk25) then
                pixel_data_from_rom <= image_data(address);
                pixel_pkq <= pkq(address);
          
        end if;
           
    end process;
end Behavioral;
